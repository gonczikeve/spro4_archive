----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/11/2023 01:08:29 AM
-- Design Name: 
-- Module Name: filter_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;
--use IEEE.std_logic_arith.all;
--use ieee.std_logic_unsigned.all;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity filter2_tb is
--  Port ( );
end filter2_tb;

architecture Behavioral2 of filter2_tb is
    component sine_signed is
        Port (wave_out: out std_logic_vector(23 downto 0);
    clock: in std_logic;
    reset: in std_logic);
    end component;
    
    component filter2 is
    Port ( Clock : in STD_LOGIC;
           Data : in STD_LOGIC_VECTOR (23 downto 0);
           data_out : out  STD_LOGIC_VECTOR(23 downto 0);
           reset : in STD_LOGIC;
           coefficients: in std_logic_vector(3719 downto 0));
    end component;
    
    
    signal Clock: std_logic;
    signal clockdiv: std_logic :='0';
    signal sin_to_filter: std_logic_vector(23 downto 0);
    --signal sin1_out: std_logic_vector(15 downto 0);
    signal sin2_out: STD_LOGIC_VECTOR(23 downto 0);
    --signal sinadder: std_logic_vector(15 downto 0);
    --signal toadder1:std_logic_vector(15 downto 0);
    --signal toadder2:std_logic_vector(15 downto 0);
    
begin
    --sinadder <= toadder1 + toadder2;
    
    sine_gen: sine_signed port map(Clock => Clock, wave_out => sin_to_filter, reset => '0');
    --sine_gen2: sine port map(Clock => clockdiv, result => toadder2);
    filterUT: filter2 port map(Clock => Clock, Data => sin_to_filter, data_out => sin2_out, reset=> '0', coefficients =>
   "000000000000000010001010000000000000001110011110000000000000011010010011000000000000100100111010000000000000101101100110000000000000110011100011000000000000110101111111000000000000110100001101000000000000101101101011000000000000100010000110000000000000010001100011011001010000000000000000011010001010000000000000010110010101000000000000110111000011100000000000111010010110100000000000101110100100100000000000011011000000100000000000101011010000100000000000011000100010100000000000111010001101100000000000110100001011000000000000000000000000000110110101000000000001000001001001000000000001111110110000000000000010111010010001000000000011101101101010000000000100010010110010000000000100100011111110000000000100011100101010000000000011111001111110000000000010111011010000000000000001100010011100001100001100000000000000101011111011110000000000111111011011111000000000110111001111101000000000000011101010001000000000010110101100111100000000001110011101011100000000101111000000111100000000110001100100001000000000010110000100011000000000100111000111010000000000000000000000010001010100000000000100000011001100000000000111111100000010000000001011100110100100000000001110101100001001000000010000110110101110000000010001110010101101000000010001010001000001000000001111001000110011000000001011011000111101000000000110001001000010001101100110000000000000111010001010001000000000010100010101000100000000100010010010100110000000111001111011010010000000110000011000011111000000100110111001110111000000011100000000001111000000110111001101111111000000010100111111011010000000010011110111100100000000000000000000011001101111000000010010000001101000000000100110001110011011000000111100001111000010000001010011001000101110000001101001111010010111000001111111100000001001000010010010110111100000000010100011000011010010000010101111001111011001000010110110110100000110000010111001011000011111000010110110110100000110000010101111001111011001000010100011000011010010000010010010110111100000000001111111100000001001000001101001111010010111000001010011001000101110000000111100001111000010000000100110001110011011000000010010000001101000000000000000011001101111010011110111100100000000010100111111011010000000110111001101111111000000011100000000001111000000100110111001110111000000110000011000011111000000111001111011010010000000100010010010100110000000010100010101000100000000111010001010001000000000001101100110000000000000000000000110001001000010000000001011011000111101000000001111001000110011000000010001010001000001000000010001110010101101000000010000110110101110000000001110101100001001000000001011100110100100000000000111111100000010000000000100000011001100000000000000010001010100100111000111010000000000010110000100011000000000110001100100001000000000101111000000111100000000001110011101011100000000010110101100111100000000000011101010001000000000110111001111101000000000111111011011111000000000101011111011110000000000001100001100000000000000000000000001100010011100000000000010111011010000000000000011111001111110000000000100011100101010000000000100100011111110000000000100010010110010000000000011101101101010000000000010111010010001000000000001111110110000000000000001000001001001000000000000000110110101110100001011000000000000111010001101100000000000011000100010100000000000101011010000100000000000011011000000100000000000101110100100100000000000111010010110100000000000110111000011100000000000010110010101000000000000011010001010000000000000011001010000000000000000000000000000010001100011000000000000100010000110000000000000101101101011000000000000110100001101000000000000110101111111000000000000110011100011000000000000101101100110000000000000100100111010000000000000011010010011000000000000001110011110000000000000000010001010");                  
    Clock_process: process
    begin
        clock <= '0';
        clockdiv <= not clockdiv;
        wait for 11338 ns;
        clock <= '1';
        wait for 11338 ns;
    end process;
end Behavioral2;
