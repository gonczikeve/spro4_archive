----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 04/30/2023 01:54:28 PM
-- Design Name: 
-- Module Name: sine_signed - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity sine_signed is
    Port (
    clock: in std_logic;
    wave_out: out std_logic_vector(23 downto 0):=(others =>'0');
    reset: in std_logic);
end sine_signed;

architecture Behavioral3 of sine_signed is

type table_type is array(0 to 440) of integer;
    constant sin_table: table_type := (
        0, 119513, 239002, 358443, 477811, 597082, 716231, 835236, 954070, 1072711, 
1191135, 1309316, 1427232, 1544858, 1662170, 1779145, 1895759, 2011988, 2127809, 2243197, 
2358131, 2472585, 2586538, 2699966, 2812845, 2925154, 3036869, 3147967, 3258427, 3368225, 
3477339, 3585748, 3693428, 3800359, 3906518, 4011885, 4116437, 4220153, 4323013, 4424995, 
4526079, 4626244, 4725471, 4823738, 4921025, 5017314, 5112585, 5206817, 5299993, 5392093, 
5483098, 5572990, 5661751, 5749363, 5835808, 5921068, 6005126, 6087965, 6169568, 6249919, 
6329001, 6406799, 6483296, 6558477, 6632327, 6704830, 6775973, 6845739, 6914117, 6981091, 
7046647, 7110774, 7173457, 7234683, 7294442, 7352719, 7409504, 7464785, 7518551, 7570790, 
7621493, 7670648, 7718247, 7764278, 7808734, 7851605, 7892881, 7932556, 7970620, 8007067, 
8041888, 8075076, 8106626, 8136530, 8164782, 8191377, 8216309, 8239573, 8261165, 8281080, 
8299314, 8315863, 8330724, 8343894, 8355370, 8365151, 8373233, 8379616, 8384297, 8387277, 
8388554, 8388128, 8386000, 8382169, 8376637, 8369404, 8360473, 8349844, 8337521, 8323505, 
8307799, 8290407, 8271332, 8250579, 8228150, 8204051, 8178287, 8150863, 8121784, 8091057, 
8058687, 8024681, 7989046, 7951790, 7912919, 7872443, 7830368, 7786704, 7741459, 7694643, 
7646264, 7596334, 7544862, 7491858, 7437333, 7381299, 7323766, 7264747, 7204253, 7142296, 
7078890, 7014047, 6947780, 6880103, 6811029, 6740572, 6668748, 6595569, 6521052, 6445211, 
6368062, 6289620, 6209901, 6128922, 6046699, 5963248, 5878587, 5792732, 5705702, 5617513, 
5528184, 5437733, 5346178, 5253538, 5159832, 5065078, 4969296, 4872505, 4774725, 4675976, 
4576278, 4475651, 4374115, 4271691, 4168401, 4064264, 3959302, 3853536, 3746989, 3639680, 
3531633, 3422869, 3313410, 3203278, 3092497, 2981087, 2869073, 2756476, 2643319, 2529626, 
2415419, 2300722, 2185558, 2069951, 1953923, 1837499, 1720701, 1603555, 1486082, 1368309, 
1250257, 1131952, 1013416, 894676, 775753, 656673, 537460, 418138, 298730, 179262, 
59758, -59758, -179262, -298730, -418138, -537460, -656673, -775753, -894676, -1013416, 
-1131952, -1250257, -1368309, -1486082, -1603555, -1720701, -1837499, -1953923, -2069951, -2185558, 
-2300722, -2415419, -2529626, -2643319, -2756476, -2869073, -2981087, -3092497, -3203278, -3313410, 
-3422869, -3531633, -3639680, -3746989, -3853536, -3959302, -4064264, -4168401, -4271691, -4374115, 
-4475651, -4576278, -4675976, -4774725, -4872505, -4969296, -5065078, -5159832, -5253538, -5346178, 
-5437733, -5528184, -5617513, -5705702, -5792732, -5878587, -5963248, -6046699, -6128922, -6209901, 
-6289620, -6368062, -6445211, -6521052, -6595569, -6668748, -6740572, -6811029, -6880103, -6947780, 
-7014047, -7078890, -7142296, -7204253, -7264747, -7323766, -7381299, -7437333, -7491858, -7544862, 
-7596334, -7646264, -7694643, -7741459, -7786704, -7830368, -7872443, -7912919, -7951790, -7989046, 
-8024681, -8058687, -8091057, -8121784, -8150863, -8178287, -8204051, -8228150, -8250579, -8271332, 
-8290407, -8307799, -8323505, -8337521, -8349844, -8360473, -8369404, -8376637, -8382169, -8386000, 
-8388128, -8388554, -8387277, -8384297, -8379616, -8373233, -8365151, -8355370, -8343894, -8330724, 
-8315863, -8299314, -8281080, -8261165, -8239573, -8216309, -8191377, -8164782, -8136530, -8106626, 
-8075076, -8041888, -8007067, -7970620, -7932556, -7892881, -7851605, -7808734, -7764278, -7718247, 
-7670648, -7621493, -7570790, -7518551, -7464785, -7409504, -7352719, -7294442, -7234683, -7173457, 
-7110774, -7046647, -6981091, -6914117, -6845739, -6775973, -6704830, -6632327, -6558477, -6483296, 
-6406799, -6329001, -6249919, -6169568, -6087965, -6005126, -5921068, -5835808, -5749363, -5661751, 
-5572990, -5483098, -5392093, -5299993, -5206817, -5112585, -5017314, -4921025, -4823738, -4725471, 
-4626244, -4526079, -4424995, -4323013, -4220153, -4116437, -4011885, -3906518, -3800359, -3693428, 
-3585748, -3477339, -3368225, -3258427, -3147967, -3036869, -2925154, -2812845, -2699966, -2586538, 
-2472585, -2358131, -2243197, -2127809, -2011988, -1895759, -1779145, -1662170, -1544858, -1427232, 
-1309316, -1191135, -1072711, -954070, -835236, -716231, -597082, -477811, -358443, -239002, 
-119513);

begin
process(Clock)
    variable counter: integer range 0 to 441 := 0;
    variable counter2: integer range 0 to 441 :=0;
begin
    if rising_edge(clock) then
        
        wave_out <= std_logic_vector(shift_right(to_signed(sin_table(counter),24),1) + shift_right(to_signed(sin_table(counter2),24),1));
        counter := counter+1;
        counter2 := counter2+2;
        if counter = 441 then
                counter := 0;
        end if;
        if counter2 = 440 then
                counter2 := 0;
        end if;
    end if;
end process;
    
end Behavioral3;
