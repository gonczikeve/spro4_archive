----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 05/08/2023 04:15:04 PM
-- Design Name: 
-- Module Name: synth_tb - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity synth_tb is
--  Port ( );
    generic(
        coeff_bitwidth: integer:= 16;
        coeff_count: integer:=201;
        din_bitwidth: integer:=24;
        dout_bitwidth: integer:=24);
    Port (
           CLock : in STD_LOGIC;
           Data : in STD_LOGIC_VECTOR (din_bitwidth-1 downto 0);
           data_out : out STD_LOGIC_VECTOR (dout_bitwidth-1 downto 0);
           reset : in STD_LOGIC);
           --coefficients: in signed(coeff_bitwidth * coeff_count-1  downto 0));
end synth_tb;

architecture Behavioral of synth_tb is
    component filter2 is
    generic(
        coeff_bitwidth: integer:= 16;
        coeff_count: integer:=201;
        din_bitwidth: integer:=24;
        dout_bitwidth: integer:=24);
    Port ( Clock : in STD_LOGIC;
           Data : in STD_LOGIC_VECTOR (din_bitwidth-1 downto 0);
           data_out : out  STD_LOGIC_VECTOR(dout_bitwidth-1 downto 0);
           reset : in STD_LOGIC;
           coefficients: in signed(coeff_count*coeff_bitwidth-1 downto 0));
    end component;
    
    
begin
filterUT: filter2 generic map(coeff_count => coeff_count,coeff_bitwidth => coeff_bitwidth)
   port map(Clock => clock, Data => Data, data_out => data_out, reset=> '0', coefficients =>"101000000000000010100000000000001010000000000000101000000000000010100000000000001010000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000111000000000000011100000000000001110000000000000010000000000000001000000000000001100000000000000110000000000000010000000000000000000000000000000000000000000000100000000000000100000000000000011000000000000010100000000000001100000000000001000000000000000101000000000000011000000000000001110000000000001000000000000000100110000000000010110000000000001100100000000000111000000000000100000000000000010001100000000001001110000000000101011000000000011000000000000001101000000000000111001000000000011111000000000010001000000000001001001000000000100111100000000010101010000000001011011000000000110001000000000011010010000000001101111000000000111011100000000011111100000000010000101000000001000110100000000100101010000000010011101000000001010010100000000101011010000000010110110000000001011111000000000110001110000000011010000000000001101100100000000111000010000000011101010000000001111001100000000111111000000000100000101000000010000111000000001000101110000000100011111000000010010100000000001001100010000000100111001000000010100000100000001010010100000000101010001000000010101100100000001011000010000000101101000000000010110111100000001011101100000000101111101000000011000001100000001100010010000000110001111000000011001010000000001100110010000000110011101000000011010001000000001101001100000000110101001000000011010110000000001101011110000000110110001000000011011001100000001101101010000000110110110000000011011011000000001101101110000000110110110000000011011011000000001101101010000000110110011000000011011000100000001101011110000000110101100000000011010100100000001101001100000000110100010000000011001110100000001100110010000000110010100000000011000111100000001100010010000000110000011000000010111110100000001011101100000000101101111000000010110100000000001011000010000000101011001000000010101000100000001010010100000000101000001000000010011100100000001001100010000000100101000000000010001111100000001000101110000000100001110000000010000010100000000111111000000000011110011000000001110101000000000111000010000000011011001000000001101000000000000110001110000000010111110000000001011011000000000101011010000000010100101000000001001110100000000100101010000000010001101000000001000010100000000011111100000000001110111000000000110111100000000011010010000000001100010000000000101101100000000010101010000000001001111000000000100100100000000010001000000000000111110000000000011100100000000001101000000000000110000000000000010101100000000001001110000000000100011000000000010000000000000000111000000000000011001000000000001011000000000000100110000000000010000000000000000111000000000000011000000000000001010000000000000100000000000000001100000000000000101000000000000001100000000000000100000000000000001000000000000000010000000000000001100000000000000110000000000000001000000000000000100000000000000111000000000000011100000000000001110000000000000011000000000000001100000000000000110000000000000011000000000000001100000000000000110000000000000101000000000000010100000000000001010000000000000101000000000000010100000000000001010000000000000");
end Behavioral;
